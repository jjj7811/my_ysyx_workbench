//Generate the verilog at 2024-02-29T01:44:42
module top (
clk,
out,
a,
b,
op,
result
);

input clk ;
output out ;
input [3:0] a ;
input [3:0] b ;
input [2:0] op ;
output [3:0] result ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire _136_ ;
wire \op[0] ;
wire \op[2] ;
wire \op[1] ;
wire \b[0] ;
wire \b[1] ;
wire \b[2] ;
wire \b[3] ;
wire \a[3] ;
wire \a[2] ;
wire \a[1] ;
wire \a[0] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire clk ;
wire out ;

CLKBUF_X1 _137_ ( .A(_024_ ), .Z(_010_ ) );
XOR2_X2 _138_ ( .A(_024_ ), .B(_025_ ), .Z(_054_ ) );
INV_X32 _139_ ( .A(_123_ ), .ZN(_055_ ) );
NAND2_X4 _140_ ( .A1(_055_ ), .A2(_122_ ), .ZN(_056_ ) );
NOR2_X1 _141_ ( .A1(_056_ ), .A2(_124_ ), .ZN(_057_ ) );
MUX2_X1 _142_ ( .A(_025_ ), .B(_054_ ), .S(_057_ ), .Z(_011_ ) );
NOR2_X4 _143_ ( .A1(_024_ ), .A2(_025_ ), .ZN(_058_ ) );
XNOR2_X2 _144_ ( .A(_058_ ), .B(_026_ ), .ZN(_059_ ) );
MUX2_X1 _145_ ( .A(_026_ ), .B(_059_ ), .S(_057_ ), .Z(_012_ ) );
INV_X8 _146_ ( .A(_026_ ), .ZN(_060_ ) );
AND2_X2 _147_ ( .A1(_058_ ), .A2(_060_ ), .ZN(_061_ ) );
INV_X2 _148_ ( .A(_027_ ), .ZN(_062_ ) );
XNOR2_X1 _149_ ( .A(_061_ ), .B(_062_ ), .ZN(_063_ ) );
AND2_X1 _150_ ( .A1(_063_ ), .A2(_057_ ), .ZN(_064_ ) );
INV_X1 _151_ ( .A(_057_ ), .ZN(_065_ ) );
AOI21_X1 _152_ ( .A(_064_ ), .B1(_062_ ), .B2(_065_ ), .ZN(_013_ ) );
INV_X1 _153_ ( .A(_021_ ), .ZN(_066_ ) );
XNOR2_X1 _154_ ( .A(_059_ ), .B(_066_ ), .ZN(_067_ ) );
INV_X2 _155_ ( .A(_067_ ), .ZN(_068_ ) );
XNOR2_X2 _156_ ( .A(_025_ ), .B(_020_ ), .ZN(_069_ ) );
AND2_X4 _157_ ( .A1(_024_ ), .A2(_019_ ), .ZN(_070_ ) );
AND2_X4 _158_ ( .A1(_069_ ), .A2(_070_ ), .ZN(_071_ ) );
AOI21_X4 _159_ ( .A(_071_ ), .B1(_020_ ), .B2(_054_ ), .ZN(_072_ ) );
NOR2_X2 _160_ ( .A1(_068_ ), .A2(_072_ ), .ZN(_073_ ) );
AOI21_X2 _161_ ( .A(_073_ ), .B1(_021_ ), .B2(_059_ ), .ZN(_074_ ) );
INV_X1 _162_ ( .A(_022_ ), .ZN(_075_ ) );
XNOR2_X1 _163_ ( .A(_063_ ), .B(_075_ ), .ZN(_076_ ) );
NOR2_X2 _164_ ( .A1(_074_ ), .A2(_076_ ), .ZN(_077_ ) );
NOR2_X1 _165_ ( .A1(_063_ ), .A2(_075_ ), .ZN(_078_ ) );
OAI21_X1 _166_ ( .A(_057_ ), .B1(_077_ ), .B2(_078_ ), .ZN(_079_ ) );
NOR2_X1 _167_ ( .A1(_124_ ), .A2(_123_ ), .ZN(_080_ ) );
INV_X1 _168_ ( .A(_122_ ), .ZN(_081_ ) );
AND2_X1 _169_ ( .A1(_080_ ), .A2(_081_ ), .ZN(_082_ ) );
INV_X1 _170_ ( .A(_082_ ), .ZN(_083_ ) );
AOI21_X1 _171_ ( .A(_083_ ), .B1(_062_ ), .B2(_075_ ), .ZN(_084_ ) );
XNOR2_X2 _172_ ( .A(_026_ ), .B(_021_ ), .ZN(_085_ ) );
NAND2_X1 _173_ ( .A1(_025_ ), .A2(_020_ ), .ZN(_086_ ) );
OAI211_X2 _174_ ( .A(_024_ ), .B(_019_ ), .C1(_025_ ), .C2(_020_ ), .ZN(_087_ ) );
AOI21_X1 _175_ ( .A(_085_ ), .B1(_086_ ), .B2(_087_ ), .ZN(_088_ ) );
INV_X1 _176_ ( .A(_088_ ), .ZN(_089_ ) );
NAND2_X1 _177_ ( .A1(_026_ ), .A2(_021_ ), .ZN(_090_ ) );
NAND2_X1 _178_ ( .A1(_089_ ), .A2(_090_ ), .ZN(_091_ ) );
AND2_X1 _179_ ( .A1(_027_ ), .A2(_022_ ), .ZN(_092_ ) );
OAI21_X1 _180_ ( .A(_084_ ), .B1(_091_ ), .B2(_092_ ), .ZN(_093_ ) );
OAI211_X2 _181_ ( .A(_079_ ), .B(_093_ ), .C1(_023_ ), .C2(_080_ ), .ZN(_014_ ) );
XNOR2_X1 _182_ ( .A(_027_ ), .B(_022_ ), .ZN(_094_ ) );
OAI21_X1 _183_ ( .A(_094_ ), .B1(_060_ ), .B2(_021_ ), .ZN(_095_ ) );
XOR2_X2 _184_ ( .A(_024_ ), .B(_019_ ), .Z(_096_ ) );
INV_X1 _185_ ( .A(_096_ ), .ZN(_097_ ) );
AOI22_X1 _186_ ( .A1(_097_ ), .A2(_069_ ), .B1(_060_ ), .B2(_021_ ), .ZN(_098_ ) );
INV_X1 _187_ ( .A(_019_ ), .ZN(_099_ ) );
INV_X16 _188_ ( .A(_020_ ), .ZN(_100_ ) );
AOI211_X2 _189_ ( .A(_024_ ), .B(_099_ ), .C1(_025_ ), .C2(_100_ ), .ZN(_101_ ) );
NOR2_X1 _190_ ( .A1(_100_ ), .A2(_025_ ), .ZN(_102_ ) );
NOR2_X1 _191_ ( .A1(_101_ ), .A2(_102_ ), .ZN(_103_ ) );
AOI21_X1 _192_ ( .A(_095_ ), .B1(_098_ ), .B2(_103_ ), .ZN(_104_ ) );
INV_X16 _193_ ( .A(_124_ ), .ZN(_105_ ) );
NOR2_X2 _194_ ( .A1(_105_ ), .A2(_122_ ), .ZN(_106_ ) );
OAI211_X2 _195_ ( .A(_106_ ), .B(_123_ ), .C1(_062_ ), .C2(_022_ ), .ZN(_107_ ) );
OR2_X2 _196_ ( .A1(_104_ ), .A2(_107_ ), .ZN(_108_ ) );
AND2_X1 _197_ ( .A1(_122_ ), .A2(_123_ ), .ZN(_109_ ) );
AND4_X1 _198_ ( .A1(_124_ ), .A2(_085_ ), .A3(_094_ ), .A4(_109_ ), .ZN(_110_ ) );
NAND3_X1 _199_ ( .A1(_110_ ), .A2(_069_ ), .A3(_097_ ), .ZN(_111_ ) );
OAI211_X2 _200_ ( .A(_106_ ), .B(_055_ ), .C1(_024_ ), .C2(_019_ ), .ZN(_112_ ) );
NAND4_X1 _201_ ( .A1(_096_ ), .A2(_122_ ), .A3(_124_ ), .A4(_055_ ), .ZN(_113_ ) );
AND4_X2 _202_ ( .A1(_108_ ), .A2(_111_ ), .A3(_112_ ), .A4(_113_ ), .ZN(_114_ ) );
BUF_X4 _203_ ( .A(_105_ ), .Z(_115_ ) );
AND3_X1 _204_ ( .A1(_109_ ), .A2(_070_ ), .A3(_115_ ), .ZN(_116_ ) );
NOR2_X1 _205_ ( .A1(_055_ ), .A2(_122_ ), .ZN(_117_ ) );
AND2_X1 _206_ ( .A1(_117_ ), .A2(_115_ ), .ZN(_118_ ) );
AOI221_X4 _207_ ( .A(_116_ ), .B1(_096_ ), .B2(_057_ ), .C1(_099_ ), .C2(_118_ ), .ZN(_119_ ) );
OAI211_X2 _208_ ( .A(_114_ ), .B(_119_ ), .C1(_083_ ), .C2(_097_ ), .ZN(_015_ ) );
AOI211_X4 _209_ ( .A(_124_ ), .B(_056_ ), .C1(_069_ ), .C2(_070_ ), .ZN(_120_ ) );
XNOR2_X1 _210_ ( .A(_054_ ), .B(_100_ ), .ZN(_121_ ) );
OAI21_X1 _211_ ( .A(_120_ ), .B1(_121_ ), .B2(_070_ ), .ZN(_028_ ) );
NOR2_X1 _212_ ( .A1(_069_ ), .A2(_070_ ), .ZN(_029_ ) );
OAI21_X1 _213_ ( .A(_082_ ), .B1(_071_ ), .B2(_029_ ), .ZN(_030_ ) );
NAND3_X1 _214_ ( .A1(_117_ ), .A2(_115_ ), .A3(_100_ ), .ZN(_031_ ) );
NOR3_X1 _215_ ( .A1(_069_ ), .A2(_115_ ), .A3(_056_ ), .ZN(_032_ ) );
NOR2_X1 _216_ ( .A1(_025_ ), .A2(_020_ ), .ZN(_033_ ) );
NOR4_X1 _217_ ( .A1(_033_ ), .A2(_115_ ), .A3(_122_ ), .A4(_123_ ), .ZN(_034_ ) );
NAND2_X1 _218_ ( .A1(_109_ ), .A2(_115_ ), .ZN(_035_ ) );
NOR2_X1 _219_ ( .A1(_035_ ), .A2(_086_ ), .ZN(_036_ ) );
NOR3_X1 _220_ ( .A1(_032_ ), .A2(_034_ ), .A3(_036_ ), .ZN(_037_ ) );
NAND4_X1 _221_ ( .A1(_028_ ), .A2(_030_ ), .A3(_031_ ), .A4(_037_ ), .ZN(_016_ ) );
OAI21_X1 _222_ ( .A(_057_ ), .B1(_068_ ), .B2(_072_ ), .ZN(_038_ ) );
AOI21_X1 _223_ ( .A(_038_ ), .B1(_072_ ), .B2(_068_ ), .ZN(_039_ ) );
AND3_X1 _224_ ( .A1(_085_ ), .A2(_086_ ), .A3(_087_ ), .ZN(_040_ ) );
NOR3_X1 _225_ ( .A1(_040_ ), .A2(_088_ ), .A3(_083_ ), .ZN(_041_ ) );
AND3_X1 _226_ ( .A1(_117_ ), .A2(_115_ ), .A3(_066_ ), .ZN(_042_ ) );
OR3_X1 _227_ ( .A1(_085_ ), .A2(_115_ ), .A3(_056_ ), .ZN(_043_ ) );
OAI211_X2 _228_ ( .A(_106_ ), .B(_055_ ), .C1(_026_ ), .C2(_021_ ), .ZN(_044_ ) );
OAI211_X2 _229_ ( .A(_043_ ), .B(_044_ ), .C1(_035_ ), .C2(_090_ ), .ZN(_045_ ) );
OR4_X1 _230_ ( .A1(_039_ ), .A2(_041_ ), .A3(_042_ ), .A4(_045_ ), .ZN(_017_ ) );
AND3_X1 _231_ ( .A1(_109_ ), .A2(_092_ ), .A3(_115_ ), .ZN(_046_ ) );
AND2_X2 _232_ ( .A1(_074_ ), .A2(_076_ ), .ZN(_047_ ) );
NOR3_X2 _233_ ( .A1(_047_ ), .A2(_077_ ), .A3(_065_ ), .ZN(_048_ ) );
AOI211_X2 _234_ ( .A(_046_ ), .B(_048_ ), .C1(_075_ ), .C2(_118_ ), .ZN(_049_ ) );
XNOR2_X1 _235_ ( .A(_091_ ), .B(_094_ ), .ZN(_050_ ) );
NAND2_X1 _236_ ( .A1(_050_ ), .A2(_082_ ), .ZN(_051_ ) );
OAI211_X2 _237_ ( .A(_106_ ), .B(_055_ ), .C1(_027_ ), .C2(_022_ ), .ZN(_052_ ) );
OR3_X1 _238_ ( .A1(_094_ ), .A2(_115_ ), .A3(_056_ ), .ZN(_053_ ) );
NAND4_X1 _239_ ( .A1(_049_ ), .A2(_051_ ), .A3(_052_ ), .A4(_053_ ), .ZN(_018_ ) );
BUF_X1 _240_ ( .A(\op[0] ), .Z(_122_ ) );
BUF_X1 _241_ ( .A(\op[2] ), .Z(_124_ ) );
BUF_X1 _242_ ( .A(\op[1] ), .Z(_123_ ) );
BUF_X1 _243_ ( .A(\b[0] ), .Z(_024_ ) );
BUF_X1 _244_ ( .A(_010_ ), .Z(_000_ ) );
BUF_X1 _245_ ( .A(\b[1] ), .Z(_025_ ) );
BUF_X1 _246_ ( .A(_011_ ), .Z(_001_ ) );
BUF_X1 _247_ ( .A(\b[2] ), .Z(_026_ ) );
BUF_X1 _248_ ( .A(_012_ ), .Z(_002_ ) );
BUF_X1 _249_ ( .A(\b[3] ), .Z(_027_ ) );
BUF_X1 _250_ ( .A(_013_ ), .Z(_003_ ) );
BUF_X1 _251_ ( .A(\a[3] ), .Z(_022_ ) );
BUF_X1 _252_ ( .A(\a[2] ), .Z(_021_ ) );
BUF_X1 _253_ ( .A(\a[1] ), .Z(_020_ ) );
BUF_X1 _254_ ( .A(\a[0] ), .Z(_019_ ) );
BUF_X1 _255_ ( .A(_009_ ), .Z(_023_ ) );
BUF_X1 _256_ ( .A(_014_ ), .Z(_004_ ) );
BUF_X1 _257_ ( .A(\result[0] ), .Z(_125_ ) );
BUF_X1 _258_ ( .A(_015_ ), .Z(_005_ ) );
BUF_X1 _259_ ( .A(\result[1] ), .Z(_126_ ) );
BUF_X1 _260_ ( .A(_016_ ), .Z(_006_ ) );
BUF_X1 _261_ ( .A(\result[2] ), .Z(_127_ ) );
BUF_X1 _262_ ( .A(_017_ ), .Z(_007_ ) );
BUF_X1 _263_ ( .A(\result[3] ), .Z(_128_ ) );
BUF_X1 _264_ ( .A(_018_ ), .Z(_008_ ) );
DFF_X1 _265_ ( .CK(clk ), .D(_000_ ), .Q(\b[0] ), .QN(_129_ ) );
DFF_X1 _266_ ( .CK(clk ), .D(_001_ ), .Q(\b[1] ), .QN(_130_ ) );
DFF_X1 _267_ ( .CK(clk ), .D(_002_ ), .Q(\b[2] ), .QN(_131_ ) );
DFF_X1 _268_ ( .CK(clk ), .D(_003_ ), .Q(\b[3] ), .QN(_132_ ) );
DFF_X1 _269_ ( .CK(clk ), .D(_005_ ), .Q(\result[0] ), .QN(_133_ ) );
DFF_X1 _270_ ( .CK(clk ), .D(_006_ ), .Q(\result[1] ), .QN(_134_ ) );
DFF_X1 _271_ ( .CK(clk ), .D(_007_ ), .Q(\result[2] ), .QN(_135_ ) );
DFF_X1 _272_ ( .CK(clk ), .D(_008_ ), .Q(\result[3] ), .QN(_136_ ) );
DFF_X1 _273_ ( .CK(clk ), .D(_004_ ), .Q(out ), .QN(_009_ ) );

endmodule
